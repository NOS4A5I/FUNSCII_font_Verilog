/******************************************************************************
Two-color FUNSCII font bitmap.

FUNSCII font (released under CC0 license):
	https://github.com/Wuerfel21/funscii/blob/master/LICENSE-font.txt

The original memory source (font.bin) found here:
	https://forums.parallax.com/discussion/167894/a-rom-font-compatible-8x8-font
******************************************************************************/

// FUNSCII Font ROM module
//
// Input:
//
//      [7:0] char_idx : A character index, ranging 0-255.
//
// Output:
//
//      [0:63] char_out : The 8x8 bitmap output of the character
//      at that index. First 8 bits [0:7] are the first row of the 8x8 character,
//      next 8 bits [8:15] are the next row, etc.
//
module funscii_font(
    input [7:0] char_idx, // up to 256 accessible characters
    output reg [0:63] char_out // 64 pixels out (8x8 bitmap)
);

    reg [0:16383] font_mem = {
        8'hFF, 8'h80, 8'hB0, 8'hA0, 8'hA0, 8'hB0, 8'h80, 8'h80, 8'hFF, 8'h80, 8'h80, 8'h80,
        8'h80, 8'h80, 8'h80, 8'hFF, 8'h00, 8'h10, 8'h30, 8'h7F, 8'h7F, 8'h30, 8'h10, 8'h00,
        8'h00, 8'h08, 8'h0C, 8'hFE, 8'hFE, 8'h0C, 8'h08, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18,
        8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18,
        8'h03, 8'h0F, 8'h3F, 8'hFF, 8'h3F, 8'h0F, 8'h03, 8'h00, 8'hC0, 8'hF0, 8'hFC, 8'hFF,
        8'hFC, 8'hF0, 8'hC0, 8'h00, 8'hFF, 8'h00, 8'h06, 8'h02, 8'h02, 8'h06, 8'h00, 8'h00,
        8'hFF, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'hFF, 8'h80, 8'h80, 8'h80, 8'h80,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'h80, 8'h80, 8'h01, 8'h01, 8'h01, 8'h01,
        8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00,
        8'h00, 8'h00, 8'h00, 8'hFF, 8'h3C, 8'h7E, 8'h7E, 8'h7E, 8'h7E, 8'h7E, 8'h3C, 8'h00,
        8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6,
        8'hC6, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'hFE, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h00,
        8'hFE, 8'h60, 8'h30, 8'h18, 8'h30, 8'h60, 8'hFE, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6,
        8'hC6, 8'h6C, 8'hEE, 8'h00, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h00,
        8'h01, 8'h03, 8'h06, 8'h8C, 8'hD8, 8'h70, 8'h20, 8'h00, 8'h06, 8'h0E, 8'h76, 8'h06,
        8'h06, 8'h00, 8'h00, 8'h00, 8'h02, 8'h04, 8'h08, 8'h10, 8'h30, 8'h50, 8'h90, 8'h10,
        8'h10, 8'h10, 8'h10, 8'hFE, 8'h82, 8'h44, 8'h28, 8'h10, 8'h09, 8'h09, 8'h09, 8'hF9,
        8'h09, 8'h09, 8'h09, 8'h00, 8'h09, 8'h09, 8'h69, 8'h99, 8'h69, 8'h09, 8'h09, 8'h00,
        8'h10, 8'hF0, 8'h00, 8'h00, 8'h00, 8'hF0, 8'h10, 8'h10, 8'h01, 8'h01, 8'h01, 8'hFF,
        8'h01, 8'h01, 8'h01, 8'h00, 8'h01, 8'h31, 8'h19, 8'h01, 8'h31, 8'h19, 8'h01, 8'h00,
        8'h10, 8'h20, 8'h40, 8'h80, 8'h90, 8'h50, 8'h30, 8'hF0, 8'h90, 8'hA0, 8'hC0, 8'hF0,
        8'h80, 8'h40, 8'h20, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
        8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h00, 8'h66, 8'h66, 8'h66, 8'h00,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h6C, 8'h6C, 8'hFE, 8'h6C, 8'hFE, 8'h6C, 8'h6C, 8'h00,
        8'h18, 8'h3E, 8'h60, 8'h3C, 8'h06, 8'h7C, 8'h18, 8'h00, 8'h00, 8'hC6, 8'hCC, 8'h18,
        8'h30, 8'h66, 8'hC6, 8'h00, 8'h38, 8'h6C, 8'h38, 8'h76, 8'hDC, 8'hCC, 8'h76, 8'h00,
        8'h18, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h18, 8'h30, 8'h30,
        8'h30, 8'h18, 8'h0C, 8'h00, 8'h30, 8'h18, 8'h0C, 8'h0C, 8'h0C, 8'h18, 8'h30, 8'h00,
        8'h00, 8'h66, 8'h3C, 8'hFF, 8'h3C, 8'h66, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h7E,
        8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h30,
        8'h00, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
        8'h00, 8'h18, 8'h18, 8'h00, 8'h03, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'h00,
        8'h3C, 8'h66, 8'h6E, 8'h76, 8'h66, 8'h66, 8'h3C, 8'h00, 8'h18, 8'h38, 8'h18, 8'h18,
        8'h18, 8'h18, 8'h7E, 8'h00, 8'h3C, 8'h66, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h7E, 8'h00,
        8'h3C, 8'h66, 8'h06, 8'h1C, 8'h06, 8'h66, 8'h3C, 8'h00, 8'h1C, 8'h3C, 8'h6C, 8'hCC,
        8'hFE, 8'h0C, 8'h0C, 8'h00, 8'h7E, 8'h60, 8'h7C, 8'h06, 8'h06, 8'h66, 8'h3C, 8'h00,
        8'h1C, 8'h30, 8'h60, 8'h7C, 8'h66, 8'h66, 8'h3C, 8'h00, 8'h7E, 8'h06, 8'h06, 8'h0C,
        8'h18, 8'h18, 8'h18, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h3C, 8'h66, 8'h66, 8'h3C, 8'h00,
        8'h3C, 8'h66, 8'h66, 8'h3E, 8'h06, 8'h0C, 8'h38, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00,
        8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h18, 8'h18, 8'h30,
        8'h0C, 8'h18, 8'h30, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h00,
        8'h7E, 8'h00, 8'h00, 8'h00, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h00,
        8'h3C, 8'h66, 8'h06, 8'h0C, 8'h18, 8'h00, 8'h18, 8'h00, 8'h7C, 8'hC6, 8'hDE, 8'hDE,
        8'hDE, 8'hC0, 8'h7C, 8'h00, 8'h18, 8'h3C, 8'h66, 8'h66, 8'h7E, 8'h66, 8'h66, 8'h00,
        8'h7C, 8'h66, 8'h66, 8'h7C, 8'h66, 8'h66, 8'h7C, 8'h00, 8'h3C, 8'h66, 8'h60, 8'h60,
        8'h60, 8'h66, 8'h3C, 8'h00, 8'h78, 8'h6C, 8'h66, 8'h66, 8'h66, 8'h6C, 8'h78, 8'h00,
        8'h7E, 8'h60, 8'h60, 8'h7C, 8'h60, 8'h60, 8'h7E, 8'h00, 8'h7E, 8'h60, 8'h60, 8'h7C,
        8'h60, 8'h60, 8'h60, 8'h00, 8'h3C, 8'h66, 8'h60, 8'h6E, 8'h66, 8'h66, 8'h3E, 8'h00,
        8'h66, 8'h66, 8'h66, 8'h7E, 8'h66, 8'h66, 8'h66, 8'h00, 8'h7E, 8'h18, 8'h18, 8'h18,
        8'h18, 8'h18, 8'h7E, 8'h00, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h66, 8'h3C, 8'h00,
        8'hC6, 8'hCC, 8'hD8, 8'hF0, 8'hD8, 8'hCC, 8'hC6, 8'h00, 8'h60, 8'h60, 8'h60, 8'h60,
        8'h60, 8'h60, 8'h7E, 8'h00, 8'hC6, 8'hEE, 8'hFE, 8'hD6, 8'hC6, 8'hC6, 8'hC6, 8'h00,
        8'hC6, 8'hE6, 8'hF6, 8'hDE, 8'hCE, 8'hC6, 8'hC6, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66,
        8'h66, 8'h66, 8'h3C, 8'h00, 8'h7C, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60, 8'h60, 8'h00,
        8'h3C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h6C, 8'h36, 8'h00, 8'h7C, 8'h66, 8'h66, 8'h7C,
        8'h6C, 8'h66, 8'h66, 8'h00, 8'h3C, 8'h66, 8'h60, 8'h3C, 8'h06, 8'h66, 8'h3C, 8'h00,
        8'h7E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66,
        8'h66, 8'h66, 8'h3C, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h18, 8'h00,
        8'hC6, 8'hC6, 8'hC6, 8'hD6, 8'hFE, 8'hEE, 8'hC6, 8'h00, 8'hC3, 8'h66, 8'h3C, 8'h18,
        8'h3C, 8'h66, 8'hC3, 8'h00, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00,
        8'h7E, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h7E, 8'h00, 8'h3C, 8'h30, 8'h30, 8'h30,
        8'h30, 8'h30, 8'h3C, 8'h00, 8'hC0, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h06, 8'h03, 8'h00,
        8'h3C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h3C, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF,
        8'h18, 8'h0C, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h06,
        8'h3E, 8'h66, 8'h3E, 8'h00, 8'h60, 8'h60, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h00,
        8'h00, 8'h00, 8'h3C, 8'h60, 8'h60, 8'h60, 8'h3C, 8'h00, 8'h06, 8'h06, 8'h3E, 8'h66,
        8'h66, 8'h66, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h60, 8'h3C, 8'h00,
        8'h1C, 8'h30, 8'h7C, 8'h30, 8'h30, 8'h30, 8'h30, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h66,
        8'h66, 8'h3E, 8'h06, 8'h7C, 8'h60, 8'h60, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00,
        8'h18, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h1E, 8'h00, 8'h0C, 8'h00, 8'h0C, 8'h0C,
        8'h0C, 8'h0C, 8'h0C, 8'h78, 8'h60, 8'h60, 8'h66, 8'h6C, 8'h78, 8'h6C, 8'h66, 8'h00,
        8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h1E, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hFE,
        8'hD6, 8'hD6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00,
        8'h00, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h7C, 8'h66,
        8'h66, 8'h7C, 8'h60, 8'h60, 8'h00, 8'h00, 8'h3E, 8'h66, 8'h66, 8'h3E, 8'h06, 8'h06,
        8'h00, 8'h00, 8'h7C, 8'h66, 8'h60, 8'h60, 8'h60, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h60,
        8'h3C, 8'h06, 8'h7C, 8'h00, 8'h30, 8'h30, 8'h7E, 8'h30, 8'h30, 8'h30, 8'h1E, 8'h00,
        8'h00, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h66, 8'h66,
        8'h66, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'hC6, 8'hC6, 8'hD6, 8'h7C, 8'h6C, 8'h00,
        8'h00, 8'h00, 8'hC6, 8'h6C, 8'h38, 8'h6C, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h66, 8'h66,
        8'h66, 8'h3E, 8'h06, 8'h3C, 8'h00, 8'h00, 8'h7E, 8'h0C, 8'h18, 8'h30, 8'h7E, 8'h00,
        8'h0E, 8'h18, 8'h18, 8'h70, 8'h18, 8'h18, 8'h0E, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18,
        8'h18, 8'h18, 8'h18, 8'h00, 8'h70, 8'h18, 8'h18, 8'h0E, 8'h18, 8'h18, 8'h70, 8'h00,
        8'h76, 8'hDC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h81, 8'h95, 8'hA9, 8'h95,
        8'hA9, 8'h95, 8'hA9, 8'h81, 8'hC3, 8'h24, 8'h24, 8'h18, 8'h24, 8'h24, 8'hC3, 8'h00,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h07, 8'h08, 8'h08, 8'h10,
        8'h20, 8'h20, 8'hC0, 8'h00, 8'h07, 8'h08, 8'h08, 8'h10, 8'h20, 8'h20, 8'hFF, 8'h00,
        8'h00, 8'h00, 8'h00, 8'h07, 8'h08, 8'h10, 8'hE0, 8'h00, 8'hC0, 8'h20, 8'h20, 8'h10,
        8'h08, 8'h08, 8'h07, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
        8'hFF, 8'h20, 8'h20, 8'h10, 8'h08, 8'h08, 8'h07, 8'h00, 8'hE0, 8'h10, 8'h08, 8'h07,
        8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'h20, 8'h20, 8'h10, 8'h08, 8'h08, 8'hFF, 8'h00,
        8'hFF, 8'h08, 8'h08, 8'h10, 8'h20, 8'h20, 8'hC0, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00,
        8'h00, 8'h00, 8'hFF, 8'h00, 8'hE0, 8'h10, 8'h08, 8'h07, 8'h08, 8'h10, 8'hE0, 8'h00,
        8'h00, 8'h00, 8'h00, 8'hE0, 8'h10, 8'h08, 8'h07, 8'h00, 8'h07, 8'h08, 8'h10, 8'hE0,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h08, 8'h10, 8'hE0, 8'h10, 8'h08, 8'h07, 8'h00,
        8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h10, 8'h10, 8'h10,
        8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'hFF, 8'h10, 8'h10, 8'h10, 8'h10,
        8'h10, 8'h10, 8'h38, 8'hFF, 8'h38, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'hF0,
        8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h1F, 8'h10, 8'h10, 8'h10, 8'h10,
        8'h10, 8'h10, 8'h10, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF,
        8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h38, 8'hF8, 8'h38, 8'h10, 8'h10, 8'h10,
        8'h10, 8'h10, 8'h38, 8'h3F, 8'h38, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h38, 8'hFF,
        8'h38, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h38, 8'hFF, 8'h38, 8'h10, 8'h10, 8'h10,
        8'h10, 8'h10, 8'h10, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h10, 8'h10, 8'h1F,
        8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hF0, 8'h10, 8'h10, 8'h10, 8'h10,
        8'h00, 8'h00, 8'h00, 8'h1F, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h38, 8'h54, 8'h92,
        8'h10, 8'h10, 8'h10, 8'h10, 8'h18, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00,
        8'h10, 8'h10, 8'h10, 8'h10, 8'h92, 8'h54, 8'h38, 8'h10, 8'h38, 8'h6C, 8'h60, 8'hF0,
        8'h60, 8'h66, 8'hFC, 8'h00, 8'h3E, 8'h60, 8'hFC, 8'h60, 8'hF8, 8'h60, 8'h3E, 8'h00,
        8'hC3, 8'h66, 8'h3C, 8'h18, 8'h3C, 8'h18, 8'h18, 8'h00, 8'h18, 8'h16, 8'h11, 8'hF0,
        8'h11, 8'h16, 8'h18, 8'h00, 8'h20, 8'h20, 8'hA0, 8'h7F, 8'hA0, 8'h20, 8'h20, 8'h00,
        8'h25, 8'h2A, 8'hA0, 8'h7F, 8'hA0, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'hC0, 8'h3F,
        8'hC0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hFC, 8'h03, 8'h00, 8'h00, 8'h00,
        8'h42, 8'h42, 8'h42, 8'hC3, 8'h42, 8'h42, 8'h42, 8'h00, 8'h00, 8'h07, 8'h00, 8'h00,
        8'h00, 8'h07, 8'h00, 8'h00, 8'h10, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h10, 8'h10,
        8'h00, 8'hC0, 8'h00, 8'h00, 8'h00, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'hFF,
        8'h80, 8'h80, 8'h00, 8'h00, 8'h3C, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
        8'h18, 8'h18, 8'h7E, 8'h18, 8'h18, 8'h00, 8'h7E, 8'h00, 8'h70, 8'h18, 8'h30, 8'h60,
        8'h78, 8'h00, 8'h00, 8'h00, 8'h78, 8'h0C, 8'h18, 8'h0C, 8'h78, 8'h00, 8'h00, 8'h00,
        8'h00, 8'h01, 8'h01, 8'hFF, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h66, 8'h66,
        8'h66, 8'h7C, 8'h60, 8'hC0, 8'h1C, 8'h22, 8'h1C, 8'h22, 8'h1C, 8'h22, 8'h1C, 8'h20,
        8'h00, 8'h00, 8'hCE, 8'h31, 8'h4A, 8'h4A, 8'h31, 8'h00, 8'h00, 8'h00, 8'h73, 8'h8C,
        8'h52, 8'h52, 8'h8C, 8'h00, 8'h30, 8'h70, 8'h30, 8'h30, 8'h30, 8'h00, 8'h00, 8'h00,
        8'h00, 8'h20, 8'h40, 8'hFF, 8'h40, 8'h20, 8'h00, 8'h00, 8'h00, 8'h04, 8'h02, 8'hFF,
        8'h02, 8'h04, 8'h00, 8'h00, 8'h0C, 8'h10, 8'h60, 8'h10, 8'h0C, 8'h10, 8'h60, 8'h10,
        8'h00, 8'h10, 8'h28, 8'hC4, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h08, 8'h14, 8'h23,
        8'h40, 8'h80, 8'h00, 8'h00, 8'h18, 8'h00, 8'h18, 8'h30, 8'h60, 8'h66, 8'h3C, 8'h00,
        8'h70, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h66, 8'h66, 8'h00, 8'h0E, 8'h00, 8'h3C, 8'h66,
        8'h7E, 8'h66, 8'h66, 8'h00, 8'h18, 8'h66, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h66, 8'h00,
        8'h76, 8'hDC, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h66, 8'h00, 8'h66, 8'h00, 8'h3C, 8'h66,
        8'h7E, 8'h66, 8'h66, 8'h00, 8'h18, 8'h18, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h66, 8'h00,
        8'h3F, 8'h6C, 8'hCC, 8'hFE, 8'hCC, 8'hCC, 8'hCF, 8'h00, 8'h3C, 8'h66, 8'h60, 8'h60,
        8'h60, 8'h66, 8'h3C, 8'h18, 8'h70, 8'h00, 8'hFE, 8'hC0, 8'hF8, 8'hC0, 8'hFE, 8'h00,
        8'h0E, 8'h00, 8'hFE, 8'hC0, 8'hF8, 8'hC0, 8'hFE, 8'h00, 8'h18, 8'h66, 8'h00, 8'hFE,
        8'hF0, 8'hC0, 8'hFE, 8'h00, 8'h66, 8'h00, 8'hFE, 8'hC0, 8'hF8, 8'hC0, 8'hFE, 8'h00,
        8'h70, 8'h00, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h0E, 8'h00, 8'h7E, 8'h18,
        8'h18, 8'h18, 8'h7E, 8'h00, 8'h18, 8'h66, 8'h00, 8'h7E, 8'h18, 8'h18, 8'h7E, 8'h00,
        8'h66, 8'h00, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h78, 8'h6C, 8'h66, 8'hF6,
        8'h66, 8'h6C, 8'h78, 8'h00, 8'h76, 8'hDC, 8'h00, 8'hC6, 8'hF6, 8'hDE, 8'hC6, 8'h00,
        8'h70, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h0E, 8'h00, 8'h7C, 8'hC6,
        8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h18, 8'h66, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h7C, 8'h00,
        8'h76, 8'hDC, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h66, 8'h00, 8'h7C, 8'hC6,
        8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'hC6, 8'h6C, 8'h38, 8'h6C, 8'hC6, 8'h00, 8'h00,
        8'h3E, 8'h66, 8'h6E, 8'h7E, 8'h76, 8'h66, 8'h7C, 8'h00, 8'h70, 8'h00, 8'hC6, 8'hC6,
        8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h0E, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00,
        8'h18, 8'h66, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h66, 8'h00, 8'hC6, 8'hC6,
        8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h0E, 8'h00, 8'h66, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h00,
        8'hC0, 8'hC0, 8'hFC, 8'hC6, 8'hFC, 8'hC0, 8'hC0, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h6C,
        8'h66, 8'h66, 8'h6C, 8'h00, 8'h70, 8'h00, 8'h3C, 8'h06, 8'h3E, 8'h66, 8'h3E, 8'h00,
        8'h0E, 8'h00, 8'h3C, 8'h06, 8'h3E, 8'h66, 8'h3E, 8'h00, 8'h18, 8'h66, 8'h00, 8'h3E,
        8'h66, 8'hC6, 8'h7E, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h3E, 8'h66, 8'hC6, 8'h7E, 8'h00,
        8'h66, 8'h00, 8'h3C, 8'h06, 8'h3E, 8'h66, 8'h3E, 8'h00, 8'h18, 8'h18, 8'h00, 8'h3E,
        8'h66, 8'hC6, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h1B, 8'h7F, 8'hD8, 8'h77, 8'h00,
        8'h00, 8'h00, 8'h3C, 8'h60, 8'h60, 8'h60, 8'h3C, 8'h18, 8'h70, 8'h00, 8'h3C, 8'h66,
        8'h7E, 8'h60, 8'h3C, 8'h00, 8'h0E, 8'h00, 8'h3C, 8'h66, 8'h7E, 8'h60, 8'h3C, 8'h00,
        8'h18, 8'h66, 8'h00, 8'h3C, 8'h7E, 8'h60, 8'h3C, 8'h00, 8'h66, 8'h00, 8'h3C, 8'h66,
        8'h7E, 8'h60, 8'h3C, 8'h00, 8'h70, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00,
        8'h0E, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h18, 8'h66, 8'h00, 8'h38,
        8'h18, 8'h18, 8'h3C, 8'h00, 8'h66, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00,
        8'h0C, 8'h3E, 8'h0C, 8'h7C, 8'hCC, 8'hCC, 8'h78, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h7C,
        8'h66, 8'h66, 8'h66, 8'h00, 8'h70, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h00,
        8'h0E, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h00, 8'h18, 8'h66, 8'h00, 8'h3C,
        8'h66, 8'h66, 8'h3C, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h3C, 8'h00,
        8'h66, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h00, 8'h18, 8'h18, 8'h00, 8'h7E,
        8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h02, 8'h7C, 8'hCE, 8'hD6, 8'hE6, 8'h7C, 8'h80,
        8'h70, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3E, 8'h00, 8'h0E, 8'h00, 8'h66, 8'h66,
        8'h66, 8'h66, 8'h3E, 8'h00, 8'h18, 8'h66, 8'h00, 8'h66, 8'h66, 8'h66, 8'h3E, 8'h00,
        8'h66, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3E, 8'h00, 8'h0E, 8'h00, 8'h66, 8'h66,
        8'h66, 8'h3E, 8'h06, 8'h3C, 8'h60, 8'h60, 8'h7C, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60,
        8'h00, 8'h00, 8'h76, 8'hDB, 8'hDB, 8'h6E, 8'h00, 8'h00
    };

    wire [13:0] idx2addr = {char_idx, 6'd0}; 
    
    integer i;
    always @(*) begin
        for (i = 0; i < 256; i = i + 1) begin
            if(i == char_idx) begin
                char_out = font_mem[i*64+:64];
            end
        end
    end
    
endmodule

// This is the testbench I used for testing access.
/*
module tb4fontmem();

    reg [7:0] idx = 0;
    wire [0:63] memout;
    
    font_rom font_mem(
        .char_idx(idx), // up to 256 accessible characters
        .char_out(memout) // 64 pixels out (8x8 bitmap)
    );
    
    initial begin
        forever begin
            #1;
            idx <= idx + 1;
        end
    end
    
    initial begin
        #257;
        $finish;
    end

endmodule
*/